/*
 * Author: 
 * Project: Harvard Architecture Processor
 * Module: Compare and Branching Instruction
 * Script:
iverilog -o cmpBrnch cmpBrnch.v cmpBrnch-tb.v
vvp cmpBrnch
gtkwave cmpBrnch.vpd
 */
module tb_cmpBrnch;

endmodule